module Practica_2
    int puto;





endmodule 
