module Practica_2






endmodule 